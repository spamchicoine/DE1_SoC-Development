// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		output wire        acl_iface_adc_sclk,                  //               acl_iface_adc.sclk
		output wire        acl_iface_adc_cs_n,                  //                            .cs_n
		input  wire        acl_iface_adc_dout,                  //                            .dout
		output wire        acl_iface_adc_din,                   //                            .din
		inout  wire        acl_iface_av_config_SDAT,            //         acl_iface_av_config.SDAT
		output wire        acl_iface_av_config_SCLK,            //                            .SCLK
		inout  wire        acl_iface_d5m_config_I2C_SDAT,       //        acl_iface_d5m_config.I2C_SDAT
		output wire        acl_iface_d5m_config_I2C_SCLK,       //                            .I2C_SCLK
		input  wire [15:0] acl_iface_d5m_config_exposure,       //                            .exposure
		output wire [5:0]  acl_iface_led_pio_export,            //           acl_iface_led_pio.export
		input  wire [3:0]  acl_iface_pushbuttons_export,        //       acl_iface_pushbuttons.export
		output wire        acl_iface_vga_CLK,                   //               acl_iface_vga.CLK
		output wire        acl_iface_vga_HS,                    //                            .HS
		output wire        acl_iface_vga_VS,                    //                            .VS
		output wire        acl_iface_vga_BLANK,                 //                            .BLANK
		output wire        acl_iface_vga_SYNC,                  //                            .SYNC
		output wire [7:0]  acl_iface_vga_R,                     //                            .R
		output wire [7:0]  acl_iface_vga_G,                     //                            .G
		output wire [7:0]  acl_iface_vga_B,                     //                            .B
		output wire        acl_iface_vga_pll_d5m_clk_clk,       //   acl_iface_vga_pll_d5m_clk.clk
		input  wire        acl_iface_vga_pll_ref_clk_clk,       //   acl_iface_vga_pll_ref_clk.clk
		input  wire        acl_iface_vga_pll_ref_reset_reset,   // acl_iface_vga_pll_ref_reset.reset
		input  wire        acl_iface_video_in_PIXEL_CLK,        //          acl_iface_video_in.PIXEL_CLK
		input  wire        acl_iface_video_in_LINE_VALID,       //                            .LINE_VALID
		input  wire        acl_iface_video_in_FRAME_VALID,      //                            .FRAME_VALID
		input  wire        acl_iface_video_in_pixel_clk_reset,  //                            .pixel_clk_reset
		input  wire [11:0] acl_iface_video_in_PIXEL_DATA,       //                            .PIXEL_DATA
		input  wire        clk_50_clk,                          //                      clk_50.clk
		output wire        kernel_clk_clk,                      //                  kernel_clk.clk
		output wire [14:0] memory_mem_a,                        //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                       //                            .mem_ba
		output wire        memory_mem_ck,                       //                            .mem_ck
		output wire        memory_mem_ck_n,                     //                            .mem_ck_n
		output wire        memory_mem_cke,                      //                            .mem_cke
		output wire        memory_mem_cs_n,                     //                            .mem_cs_n
		output wire        memory_mem_ras_n,                    //                            .mem_ras_n
		output wire        memory_mem_cas_n,                    //                            .mem_cas_n
		output wire        memory_mem_we_n,                     //                            .mem_we_n
		output wire        memory_mem_reset_n,                  //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                       //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                      //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                    //                            .mem_dqs_n
		output wire        memory_mem_odt,                      //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                       //                            .mem_dm
		input  wire        memory_oct_rzqin,                    //                            .oct_rzqin
		output wire        peripheral_hps_io_emac1_inst_TX_CLK, //                  peripheral.hps_io_emac1_inst_TX_CLK
		output wire        peripheral_hps_io_emac1_inst_TXD0,   //                            .hps_io_emac1_inst_TXD0
		output wire        peripheral_hps_io_emac1_inst_TXD1,   //                            .hps_io_emac1_inst_TXD1
		output wire        peripheral_hps_io_emac1_inst_TXD2,   //                            .hps_io_emac1_inst_TXD2
		output wire        peripheral_hps_io_emac1_inst_TXD3,   //                            .hps_io_emac1_inst_TXD3
		input  wire        peripheral_hps_io_emac1_inst_RXD0,   //                            .hps_io_emac1_inst_RXD0
		inout  wire        peripheral_hps_io_emac1_inst_MDIO,   //                            .hps_io_emac1_inst_MDIO
		output wire        peripheral_hps_io_emac1_inst_MDC,    //                            .hps_io_emac1_inst_MDC
		input  wire        peripheral_hps_io_emac1_inst_RX_CTL, //                            .hps_io_emac1_inst_RX_CTL
		output wire        peripheral_hps_io_emac1_inst_TX_CTL, //                            .hps_io_emac1_inst_TX_CTL
		input  wire        peripheral_hps_io_emac1_inst_RX_CLK, //                            .hps_io_emac1_inst_RX_CLK
		input  wire        peripheral_hps_io_emac1_inst_RXD1,   //                            .hps_io_emac1_inst_RXD1
		input  wire        peripheral_hps_io_emac1_inst_RXD2,   //                            .hps_io_emac1_inst_RXD2
		input  wire        peripheral_hps_io_emac1_inst_RXD3,   //                            .hps_io_emac1_inst_RXD3
		inout  wire        peripheral_hps_io_sdio_inst_CMD,     //                            .hps_io_sdio_inst_CMD
		inout  wire        peripheral_hps_io_sdio_inst_D0,      //                            .hps_io_sdio_inst_D0
		inout  wire        peripheral_hps_io_sdio_inst_D1,      //                            .hps_io_sdio_inst_D1
		output wire        peripheral_hps_io_sdio_inst_CLK,     //                            .hps_io_sdio_inst_CLK
		inout  wire        peripheral_hps_io_sdio_inst_D2,      //                            .hps_io_sdio_inst_D2
		inout  wire        peripheral_hps_io_sdio_inst_D3,      //                            .hps_io_sdio_inst_D3
		inout  wire        peripheral_hps_io_usb1_inst_D0,      //                            .hps_io_usb1_inst_D0
		inout  wire        peripheral_hps_io_usb1_inst_D1,      //                            .hps_io_usb1_inst_D1
		inout  wire        peripheral_hps_io_usb1_inst_D2,      //                            .hps_io_usb1_inst_D2
		inout  wire        peripheral_hps_io_usb1_inst_D3,      //                            .hps_io_usb1_inst_D3
		inout  wire        peripheral_hps_io_usb1_inst_D4,      //                            .hps_io_usb1_inst_D4
		inout  wire        peripheral_hps_io_usb1_inst_D5,      //                            .hps_io_usb1_inst_D5
		inout  wire        peripheral_hps_io_usb1_inst_D6,      //                            .hps_io_usb1_inst_D6
		inout  wire        peripheral_hps_io_usb1_inst_D7,      //                            .hps_io_usb1_inst_D7
		input  wire        peripheral_hps_io_usb1_inst_CLK,     //                            .hps_io_usb1_inst_CLK
		output wire        peripheral_hps_io_usb1_inst_STP,     //                            .hps_io_usb1_inst_STP
		input  wire        peripheral_hps_io_usb1_inst_DIR,     //                            .hps_io_usb1_inst_DIR
		input  wire        peripheral_hps_io_usb1_inst_NXT,     //                            .hps_io_usb1_inst_NXT
		input  wire        peripheral_hps_io_uart0_inst_RX,     //                            .hps_io_uart0_inst_RX
		output wire        peripheral_hps_io_uart0_inst_TX,     //                            .hps_io_uart0_inst_TX
		inout  wire        peripheral_hps_io_i2c0_inst_SDA,     //                            .hps_io_i2c0_inst_SDA
		inout  wire        peripheral_hps_io_i2c0_inst_SCL,     //                            .hps_io_i2c0_inst_SCL
		inout  wire        peripheral_hps_io_gpio_inst_GPIO53,  //                            .hps_io_gpio_inst_GPIO53
		input  wire        reset_50_reset_n                     //                    reset_50.reset_n
	);

	wire  [0:0] acl_iface_kernel_irq_irq;       // irq_mapper:sender_irq -> acl_iface:kernel_irq_irq
	wire        acl_iface_kernel_clk_clk;       // acl_iface:kernel_clk_clk -> [irq_mapper:clk, rst_controller:clk]
	wire        rst_controller_reset_out_reset; // rst_controller:reset_out -> irq_mapper:reset

	system_acl_iface acl_iface (
		.acl_internal_memorg_kernel_mode         (),                                    //       acl_internal_memorg_kernel.mode
		.acl_kernel_clk_kernel_pll_locked_export (),                                    // acl_kernel_clk_kernel_pll_locked.export
		.adc_sclk                                (acl_iface_adc_sclk),                  //                              adc.sclk
		.adc_cs_n                                (acl_iface_adc_cs_n),                  //                                 .cs_n
		.adc_dout                                (acl_iface_adc_dout),                  //                                 .dout
		.adc_din                                 (acl_iface_adc_din),                   //                                 .din
		.av_config_SDAT                          (acl_iface_av_config_SDAT),            //                        av_config.SDAT
		.av_config_SCLK                          (acl_iface_av_config_SCLK),            //                                 .SCLK
		.config_clk_clk                          (clk_50_clk),                          //                       config_clk.clk
		.d5m_config_I2C_SDAT                     (acl_iface_d5m_config_I2C_SDAT),       //                       d5m_config.I2C_SDAT
		.d5m_config_I2C_SCLK                     (acl_iface_d5m_config_I2C_SCLK),       //                                 .I2C_SCLK
		.d5m_config_exposure                     (acl_iface_d5m_config_exposure),       //                                 .exposure
		.reset_n                                 (reset_50_reset_n),                    //                     global_reset.reset_n
		.kernel_clk_clk                          (acl_iface_kernel_clk_clk),            //                       kernel_clk.clk
		.kernel_clk2x_clk                        (),                                    //                     kernel_clk2x.clk
		.kernel_clk_snoop_clk                    (kernel_clk_clk),                      //                 kernel_clk_snoop.clk
		.kernel_cra_waitrequest                  (),                                    //                       kernel_cra.waitrequest
		.kernel_cra_readdata                     (),                                    //                                 .readdata
		.kernel_cra_readdatavalid                (),                                    //                                 .readdatavalid
		.kernel_cra_burstcount                   (),                                    //                                 .burstcount
		.kernel_cra_writedata                    (),                                    //                                 .writedata
		.kernel_cra_address                      (),                                    //                                 .address
		.kernel_cra_write                        (),                                    //                                 .write
		.kernel_cra_read                         (),                                    //                                 .read
		.kernel_cra_byteenable                   (),                                    //                                 .byteenable
		.kernel_cra_debugaccess                  (),                                    //                                 .debugaccess
		.kernel_irq_irq                          (acl_iface_kernel_irq_irq),            //                       kernel_irq.irq
		.kernel_mem0_waitrequest                 (),                                    //                      kernel_mem0.waitrequest
		.kernel_mem0_readdata                    (),                                    //                                 .readdata
		.kernel_mem0_readdatavalid               (),                                    //                                 .readdatavalid
		.kernel_mem0_burstcount                  (),                                    //                                 .burstcount
		.kernel_mem0_writedata                   (),                                    //                                 .writedata
		.kernel_mem0_address                     (),                                    //                                 .address
		.kernel_mem0_write                       (),                                    //                                 .write
		.kernel_mem0_read                        (),                                    //                                 .read
		.kernel_mem0_byteenable                  (),                                    //                                 .byteenable
		.kernel_mem0_debugaccess                 (),                                    //                                 .debugaccess
		.kernel_pll_refclk_clk                   (clk_50_clk),                          //                kernel_pll_refclk.clk
		.kernel_reset_reset_n                    (),                                    //                     kernel_reset.reset_n
		.led_pio_export                          (acl_iface_led_pio_export),            //                          led_pio.export
		.memory_mem_a                            (memory_mem_a),                        //                           memory.mem_a
		.memory_mem_ba                           (memory_mem_ba),                       //                                 .mem_ba
		.memory_mem_ck                           (memory_mem_ck),                       //                                 .mem_ck
		.memory_mem_ck_n                         (memory_mem_ck_n),                     //                                 .mem_ck_n
		.memory_mem_cke                          (memory_mem_cke),                      //                                 .mem_cke
		.memory_mem_cs_n                         (memory_mem_cs_n),                     //                                 .mem_cs_n
		.memory_mem_ras_n                        (memory_mem_ras_n),                    //                                 .mem_ras_n
		.memory_mem_cas_n                        (memory_mem_cas_n),                    //                                 .mem_cas_n
		.memory_mem_we_n                         (memory_mem_we_n),                     //                                 .mem_we_n
		.memory_mem_reset_n                      (memory_mem_reset_n),                  //                                 .mem_reset_n
		.memory_mem_dq                           (memory_mem_dq),                       //                                 .mem_dq
		.memory_mem_dqs                          (memory_mem_dqs),                      //                                 .mem_dqs
		.memory_mem_dqs_n                        (memory_mem_dqs_n),                    //                                 .mem_dqs_n
		.memory_mem_odt                          (memory_mem_odt),                      //                                 .mem_odt
		.memory_mem_dm                           (memory_mem_dm),                       //                                 .mem_dm
		.memory_oct_rzqin                        (memory_oct_rzqin),                    //                                 .oct_rzqin
		.peripheral_hps_io_emac1_inst_TX_CLK     (peripheral_hps_io_emac1_inst_TX_CLK), //                       peripheral.hps_io_emac1_inst_TX_CLK
		.peripheral_hps_io_emac1_inst_TXD0       (peripheral_hps_io_emac1_inst_TXD0),   //                                 .hps_io_emac1_inst_TXD0
		.peripheral_hps_io_emac1_inst_TXD1       (peripheral_hps_io_emac1_inst_TXD1),   //                                 .hps_io_emac1_inst_TXD1
		.peripheral_hps_io_emac1_inst_TXD2       (peripheral_hps_io_emac1_inst_TXD2),   //                                 .hps_io_emac1_inst_TXD2
		.peripheral_hps_io_emac1_inst_TXD3       (peripheral_hps_io_emac1_inst_TXD3),   //                                 .hps_io_emac1_inst_TXD3
		.peripheral_hps_io_emac1_inst_RXD0       (peripheral_hps_io_emac1_inst_RXD0),   //                                 .hps_io_emac1_inst_RXD0
		.peripheral_hps_io_emac1_inst_MDIO       (peripheral_hps_io_emac1_inst_MDIO),   //                                 .hps_io_emac1_inst_MDIO
		.peripheral_hps_io_emac1_inst_MDC        (peripheral_hps_io_emac1_inst_MDC),    //                                 .hps_io_emac1_inst_MDC
		.peripheral_hps_io_emac1_inst_RX_CTL     (peripheral_hps_io_emac1_inst_RX_CTL), //                                 .hps_io_emac1_inst_RX_CTL
		.peripheral_hps_io_emac1_inst_TX_CTL     (peripheral_hps_io_emac1_inst_TX_CTL), //                                 .hps_io_emac1_inst_TX_CTL
		.peripheral_hps_io_emac1_inst_RX_CLK     (peripheral_hps_io_emac1_inst_RX_CLK), //                                 .hps_io_emac1_inst_RX_CLK
		.peripheral_hps_io_emac1_inst_RXD1       (peripheral_hps_io_emac1_inst_RXD1),   //                                 .hps_io_emac1_inst_RXD1
		.peripheral_hps_io_emac1_inst_RXD2       (peripheral_hps_io_emac1_inst_RXD2),   //                                 .hps_io_emac1_inst_RXD2
		.peripheral_hps_io_emac1_inst_RXD3       (peripheral_hps_io_emac1_inst_RXD3),   //                                 .hps_io_emac1_inst_RXD3
		.peripheral_hps_io_sdio_inst_CMD         (peripheral_hps_io_sdio_inst_CMD),     //                                 .hps_io_sdio_inst_CMD
		.peripheral_hps_io_sdio_inst_D0          (peripheral_hps_io_sdio_inst_D0),      //                                 .hps_io_sdio_inst_D0
		.peripheral_hps_io_sdio_inst_D1          (peripheral_hps_io_sdio_inst_D1),      //                                 .hps_io_sdio_inst_D1
		.peripheral_hps_io_sdio_inst_CLK         (peripheral_hps_io_sdio_inst_CLK),     //                                 .hps_io_sdio_inst_CLK
		.peripheral_hps_io_sdio_inst_D2          (peripheral_hps_io_sdio_inst_D2),      //                                 .hps_io_sdio_inst_D2
		.peripheral_hps_io_sdio_inst_D3          (peripheral_hps_io_sdio_inst_D3),      //                                 .hps_io_sdio_inst_D3
		.peripheral_hps_io_usb1_inst_D0          (peripheral_hps_io_usb1_inst_D0),      //                                 .hps_io_usb1_inst_D0
		.peripheral_hps_io_usb1_inst_D1          (peripheral_hps_io_usb1_inst_D1),      //                                 .hps_io_usb1_inst_D1
		.peripheral_hps_io_usb1_inst_D2          (peripheral_hps_io_usb1_inst_D2),      //                                 .hps_io_usb1_inst_D2
		.peripheral_hps_io_usb1_inst_D3          (peripheral_hps_io_usb1_inst_D3),      //                                 .hps_io_usb1_inst_D3
		.peripheral_hps_io_usb1_inst_D4          (peripheral_hps_io_usb1_inst_D4),      //                                 .hps_io_usb1_inst_D4
		.peripheral_hps_io_usb1_inst_D5          (peripheral_hps_io_usb1_inst_D5),      //                                 .hps_io_usb1_inst_D5
		.peripheral_hps_io_usb1_inst_D6          (peripheral_hps_io_usb1_inst_D6),      //                                 .hps_io_usb1_inst_D6
		.peripheral_hps_io_usb1_inst_D7          (peripheral_hps_io_usb1_inst_D7),      //                                 .hps_io_usb1_inst_D7
		.peripheral_hps_io_usb1_inst_CLK         (peripheral_hps_io_usb1_inst_CLK),     //                                 .hps_io_usb1_inst_CLK
		.peripheral_hps_io_usb1_inst_STP         (peripheral_hps_io_usb1_inst_STP),     //                                 .hps_io_usb1_inst_STP
		.peripheral_hps_io_usb1_inst_DIR         (peripheral_hps_io_usb1_inst_DIR),     //                                 .hps_io_usb1_inst_DIR
		.peripheral_hps_io_usb1_inst_NXT         (peripheral_hps_io_usb1_inst_NXT),     //                                 .hps_io_usb1_inst_NXT
		.peripheral_hps_io_uart0_inst_RX         (peripheral_hps_io_uart0_inst_RX),     //                                 .hps_io_uart0_inst_RX
		.peripheral_hps_io_uart0_inst_TX         (peripheral_hps_io_uart0_inst_TX),     //                                 .hps_io_uart0_inst_TX
		.peripheral_hps_io_i2c0_inst_SDA         (peripheral_hps_io_i2c0_inst_SDA),     //                                 .hps_io_i2c0_inst_SDA
		.peripheral_hps_io_i2c0_inst_SCL         (peripheral_hps_io_i2c0_inst_SCL),     //                                 .hps_io_i2c0_inst_SCL
		.peripheral_hps_io_gpio_inst_GPIO53      (peripheral_hps_io_gpio_inst_GPIO53),  //                                 .hps_io_gpio_inst_GPIO53
		.pushbuttons_export                      (acl_iface_pushbuttons_export),        //                      pushbuttons.export
		.vga_CLK                                 (acl_iface_vga_CLK),                   //                              vga.CLK
		.vga_HS                                  (acl_iface_vga_HS),                    //                                 .HS
		.vga_VS                                  (acl_iface_vga_VS),                    //                                 .VS
		.vga_BLANK                               (acl_iface_vga_BLANK),                 //                                 .BLANK
		.vga_SYNC                                (acl_iface_vga_SYNC),                  //                                 .SYNC
		.vga_R                                   (acl_iface_vga_R),                     //                                 .R
		.vga_G                                   (acl_iface_vga_G),                     //                                 .G
		.vga_B                                   (acl_iface_vga_B),                     //                                 .B
		.vga_pll_d5m_clk_clk                     (acl_iface_vga_pll_d5m_clk_clk),       //                  vga_pll_d5m_clk.clk
		.vga_pll_ref_clk_clk                     (acl_iface_vga_pll_ref_clk_clk),       //                  vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset                 (acl_iface_vga_pll_ref_reset_reset),   //                vga_pll_ref_reset.reset
		.video_in_PIXEL_CLK                      (acl_iface_video_in_PIXEL_CLK),        //                         video_in.PIXEL_CLK
		.video_in_LINE_VALID                     (acl_iface_video_in_LINE_VALID),       //                                 .LINE_VALID
		.video_in_FRAME_VALID                    (acl_iface_video_in_FRAME_VALID),      //                                 .FRAME_VALID
		.video_in_pixel_clk_reset                (acl_iface_video_in_pixel_clk_reset),  //                                 .pixel_clk_reset
		.video_in_PIXEL_DATA                     (acl_iface_video_in_PIXEL_DATA)        //                                 .PIXEL_DATA
	);

	system_irq_mapper irq_mapper (
		.clk        (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (acl_iface_kernel_irq_irq)        //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_50_reset_n),              // reset_in0.reset
		.clk            (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
